module counter();

initial
begin

$display("%t", $time);

end 
endmodule:w
 
