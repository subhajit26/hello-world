 module tb();

 initial
 begin
	 $display("suman");

 end 
 endmodule
