module hello();

initial 
begin

$display ("hello_world!");

end 
endmodule
