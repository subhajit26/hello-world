module hello();

initial 
begin

$display ("hello_world!");
$display("Done");

end 
endmodule
